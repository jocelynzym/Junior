
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h7a581def;
    ram_cell[       1] = 32'h0;  // 32'h4e8652bc;
    ram_cell[       2] = 32'h0;  // 32'hbbb23399;
    ram_cell[       3] = 32'h0;  // 32'h37569c67;
    ram_cell[       4] = 32'h0;  // 32'h6da1d5ff;
    ram_cell[       5] = 32'h0;  // 32'h96c590a7;
    ram_cell[       6] = 32'h0;  // 32'haea6b5f6;
    ram_cell[       7] = 32'h0;  // 32'hee6f57c0;
    ram_cell[       8] = 32'h0;  // 32'hccf299af;
    ram_cell[       9] = 32'h0;  // 32'hcd4776ec;
    ram_cell[      10] = 32'h0;  // 32'hb8b1d83f;
    ram_cell[      11] = 32'h0;  // 32'h1e036012;
    ram_cell[      12] = 32'h0;  // 32'h57e51b89;
    ram_cell[      13] = 32'h0;  // 32'hfa43aafc;
    ram_cell[      14] = 32'h0;  // 32'h10f75b82;
    ram_cell[      15] = 32'h0;  // 32'heb217552;
    ram_cell[      16] = 32'h0;  // 32'ha610d0da;
    ram_cell[      17] = 32'h0;  // 32'he195f873;
    ram_cell[      18] = 32'h0;  // 32'hc4be3ea4;
    ram_cell[      19] = 32'h0;  // 32'h54c467f6;
    ram_cell[      20] = 32'h0;  // 32'h74a8a4e4;
    ram_cell[      21] = 32'h0;  // 32'hd06954c5;
    ram_cell[      22] = 32'h0;  // 32'h516d0929;
    ram_cell[      23] = 32'h0;  // 32'h771c5d72;
    ram_cell[      24] = 32'h0;  // 32'h5f53ee1b;
    ram_cell[      25] = 32'h0;  // 32'h8088a79c;
    ram_cell[      26] = 32'h0;  // 32'ha1d4a6c1;
    ram_cell[      27] = 32'h0;  // 32'h4f1053b6;
    ram_cell[      28] = 32'h0;  // 32'hb0521b73;
    ram_cell[      29] = 32'h0;  // 32'hd96feb47;
    ram_cell[      30] = 32'h0;  // 32'h642f065a;
    ram_cell[      31] = 32'h0;  // 32'hf1746a6b;
    ram_cell[      32] = 32'h0;  // 32'h23fb1efa;
    ram_cell[      33] = 32'h0;  // 32'he753bdc2;
    ram_cell[      34] = 32'h0;  // 32'h540140fe;
    ram_cell[      35] = 32'h0;  // 32'h2b697c96;
    ram_cell[      36] = 32'h0;  // 32'h4de22e1f;
    ram_cell[      37] = 32'h0;  // 32'hd5be83f0;
    ram_cell[      38] = 32'h0;  // 32'h885357b0;
    ram_cell[      39] = 32'h0;  // 32'hfd2b0c0f;
    ram_cell[      40] = 32'h0;  // 32'h2e156dc1;
    ram_cell[      41] = 32'h0;  // 32'h995de65d;
    ram_cell[      42] = 32'h0;  // 32'h4a168950;
    ram_cell[      43] = 32'h0;  // 32'h6e2d4cc3;
    ram_cell[      44] = 32'h0;  // 32'h2050e3a0;
    ram_cell[      45] = 32'h0;  // 32'h7d682ff4;
    ram_cell[      46] = 32'h0;  // 32'hf2366c5c;
    ram_cell[      47] = 32'h0;  // 32'h5fa2195a;
    ram_cell[      48] = 32'h0;  // 32'ha256130f;
    ram_cell[      49] = 32'h0;  // 32'h052e9afc;
    ram_cell[      50] = 32'h0;  // 32'hce1d943c;
    ram_cell[      51] = 32'h0;  // 32'h91373635;
    ram_cell[      52] = 32'h0;  // 32'h2856f71b;
    ram_cell[      53] = 32'h0;  // 32'hef773dd1;
    ram_cell[      54] = 32'h0;  // 32'h61c214d8;
    ram_cell[      55] = 32'h0;  // 32'h7a307d05;
    ram_cell[      56] = 32'h0;  // 32'h3f763666;
    ram_cell[      57] = 32'h0;  // 32'h66510f85;
    ram_cell[      58] = 32'h0;  // 32'h03795af3;
    ram_cell[      59] = 32'h0;  // 32'h97d2e48d;
    ram_cell[      60] = 32'h0;  // 32'h6a4e5608;
    ram_cell[      61] = 32'h0;  // 32'hf31c6b48;
    ram_cell[      62] = 32'h0;  // 32'h9c01b7a9;
    ram_cell[      63] = 32'h0;  // 32'h83dcfef1;
    ram_cell[      64] = 32'h0;  // 32'h5804332e;
    ram_cell[      65] = 32'h0;  // 32'hb49c148f;
    ram_cell[      66] = 32'h0;  // 32'hf1fa04fb;
    ram_cell[      67] = 32'h0;  // 32'h98fb3ef8;
    ram_cell[      68] = 32'h0;  // 32'h31934fe5;
    ram_cell[      69] = 32'h0;  // 32'h21c903b7;
    ram_cell[      70] = 32'h0;  // 32'he6ad889a;
    ram_cell[      71] = 32'h0;  // 32'h36a8329b;
    ram_cell[      72] = 32'h0;  // 32'h30b466ce;
    ram_cell[      73] = 32'h0;  // 32'h9174e5be;
    ram_cell[      74] = 32'h0;  // 32'h57a929ef;
    ram_cell[      75] = 32'h0;  // 32'h88a18a52;
    ram_cell[      76] = 32'h0;  // 32'hbeea0886;
    ram_cell[      77] = 32'h0;  // 32'h5c29c7bd;
    ram_cell[      78] = 32'h0;  // 32'ha4094ab6;
    ram_cell[      79] = 32'h0;  // 32'h062ebd6a;
    ram_cell[      80] = 32'h0;  // 32'hacec86ec;
    ram_cell[      81] = 32'h0;  // 32'h374844e4;
    ram_cell[      82] = 32'h0;  // 32'ha63a13da;
    ram_cell[      83] = 32'h0;  // 32'hcad2faf5;
    ram_cell[      84] = 32'h0;  // 32'hc892d128;
    ram_cell[      85] = 32'h0;  // 32'hb7d2217d;
    ram_cell[      86] = 32'h0;  // 32'h63137ecc;
    ram_cell[      87] = 32'h0;  // 32'h7a272ec3;
    ram_cell[      88] = 32'h0;  // 32'h471f2694;
    ram_cell[      89] = 32'h0;  // 32'h16009527;
    ram_cell[      90] = 32'h0;  // 32'hbdf0bdab;
    ram_cell[      91] = 32'h0;  // 32'h6332bdda;
    ram_cell[      92] = 32'h0;  // 32'h6025c950;
    ram_cell[      93] = 32'h0;  // 32'h1b34bf84;
    ram_cell[      94] = 32'h0;  // 32'h6e511e3c;
    ram_cell[      95] = 32'h0;  // 32'h1555ebc7;
    ram_cell[      96] = 32'h0;  // 32'hedd645a8;
    ram_cell[      97] = 32'h0;  // 32'hb8986d4b;
    ram_cell[      98] = 32'h0;  // 32'hd941066d;
    ram_cell[      99] = 32'h0;  // 32'hcb25fd60;
    ram_cell[     100] = 32'h0;  // 32'h130035ad;
    ram_cell[     101] = 32'h0;  // 32'h8e2daccc;
    ram_cell[     102] = 32'h0;  // 32'hf861e61e;
    ram_cell[     103] = 32'h0;  // 32'h9adc43ae;
    ram_cell[     104] = 32'h0;  // 32'h935d0b90;
    ram_cell[     105] = 32'h0;  // 32'heab70938;
    ram_cell[     106] = 32'h0;  // 32'hf2525d2c;
    ram_cell[     107] = 32'h0;  // 32'h7fe60a35;
    ram_cell[     108] = 32'h0;  // 32'h69f4b441;
    ram_cell[     109] = 32'h0;  // 32'hb08ce8cb;
    ram_cell[     110] = 32'h0;  // 32'he7ecd440;
    ram_cell[     111] = 32'h0;  // 32'h9f43abc8;
    ram_cell[     112] = 32'h0;  // 32'hb4f8dbfc;
    ram_cell[     113] = 32'h0;  // 32'h99333843;
    ram_cell[     114] = 32'h0;  // 32'hd330ebf5;
    ram_cell[     115] = 32'h0;  // 32'h99bbc196;
    ram_cell[     116] = 32'h0;  // 32'h862f25a6;
    ram_cell[     117] = 32'h0;  // 32'hf25eaf3a;
    ram_cell[     118] = 32'h0;  // 32'h3a514825;
    ram_cell[     119] = 32'h0;  // 32'hc2be6ef1;
    ram_cell[     120] = 32'h0;  // 32'hcf51aa88;
    ram_cell[     121] = 32'h0;  // 32'h3d2988a0;
    ram_cell[     122] = 32'h0;  // 32'h9ae51961;
    ram_cell[     123] = 32'h0;  // 32'h23183b8f;
    ram_cell[     124] = 32'h0;  // 32'h3313ff12;
    ram_cell[     125] = 32'h0;  // 32'h0b6c934d;
    ram_cell[     126] = 32'h0;  // 32'h65ebb57a;
    ram_cell[     127] = 32'h0;  // 32'h7fae242e;
    ram_cell[     128] = 32'h0;  // 32'h203c284e;
    ram_cell[     129] = 32'h0;  // 32'hd14bca26;
    ram_cell[     130] = 32'h0;  // 32'ha7dda784;
    ram_cell[     131] = 32'h0;  // 32'h77653133;
    ram_cell[     132] = 32'h0;  // 32'h67a04e4c;
    ram_cell[     133] = 32'h0;  // 32'h0e54923a;
    ram_cell[     134] = 32'h0;  // 32'hc4683614;
    ram_cell[     135] = 32'h0;  // 32'hdf27a7bc;
    ram_cell[     136] = 32'h0;  // 32'h74743f17;
    ram_cell[     137] = 32'h0;  // 32'haced5008;
    ram_cell[     138] = 32'h0;  // 32'h17f3b451;
    ram_cell[     139] = 32'h0;  // 32'h4b781d4c;
    ram_cell[     140] = 32'h0;  // 32'h23547528;
    ram_cell[     141] = 32'h0;  // 32'hbdb78aaf;
    ram_cell[     142] = 32'h0;  // 32'he04c574a;
    ram_cell[     143] = 32'h0;  // 32'hb4e9ad0b;
    ram_cell[     144] = 32'h0;  // 32'hf2519f7f;
    ram_cell[     145] = 32'h0;  // 32'h0be59eb2;
    ram_cell[     146] = 32'h0;  // 32'h1ca2de5e;
    ram_cell[     147] = 32'h0;  // 32'hcbbc868b;
    ram_cell[     148] = 32'h0;  // 32'h7b67b4fb;
    ram_cell[     149] = 32'h0;  // 32'h22a69f13;
    ram_cell[     150] = 32'h0;  // 32'h70409687;
    ram_cell[     151] = 32'h0;  // 32'h49f93092;
    ram_cell[     152] = 32'h0;  // 32'hf42f0f43;
    ram_cell[     153] = 32'h0;  // 32'h6ea14359;
    ram_cell[     154] = 32'h0;  // 32'hdd4f4fe5;
    ram_cell[     155] = 32'h0;  // 32'hf504d4ca;
    ram_cell[     156] = 32'h0;  // 32'habd9d0de;
    ram_cell[     157] = 32'h0;  // 32'hb6a4c182;
    ram_cell[     158] = 32'h0;  // 32'hb86544a6;
    ram_cell[     159] = 32'h0;  // 32'h43ff9a0a;
    ram_cell[     160] = 32'h0;  // 32'h76b1898c;
    ram_cell[     161] = 32'h0;  // 32'h8cf3ecef;
    ram_cell[     162] = 32'h0;  // 32'h46ed7205;
    ram_cell[     163] = 32'h0;  // 32'h7343b0f6;
    ram_cell[     164] = 32'h0;  // 32'h6eb5aba2;
    ram_cell[     165] = 32'h0;  // 32'hbd648969;
    ram_cell[     166] = 32'h0;  // 32'hc1c3f766;
    ram_cell[     167] = 32'h0;  // 32'h4e9103b5;
    ram_cell[     168] = 32'h0;  // 32'hd466020e;
    ram_cell[     169] = 32'h0;  // 32'h05fa877c;
    ram_cell[     170] = 32'h0;  // 32'h0410a8e0;
    ram_cell[     171] = 32'h0;  // 32'h852f04e8;
    ram_cell[     172] = 32'h0;  // 32'ha8ddb198;
    ram_cell[     173] = 32'h0;  // 32'h8b3f63a5;
    ram_cell[     174] = 32'h0;  // 32'h2347f3bf;
    ram_cell[     175] = 32'h0;  // 32'hfdbdef06;
    ram_cell[     176] = 32'h0;  // 32'h797811cc;
    ram_cell[     177] = 32'h0;  // 32'h36cc12f9;
    ram_cell[     178] = 32'h0;  // 32'h4ef33396;
    ram_cell[     179] = 32'h0;  // 32'h4f94954a;
    ram_cell[     180] = 32'h0;  // 32'hbafe3ec0;
    ram_cell[     181] = 32'h0;  // 32'h3b7145b0;
    ram_cell[     182] = 32'h0;  // 32'h72c7c872;
    ram_cell[     183] = 32'h0;  // 32'ha889f3af;
    ram_cell[     184] = 32'h0;  // 32'hb5393ed3;
    ram_cell[     185] = 32'h0;  // 32'h19f955e9;
    ram_cell[     186] = 32'h0;  // 32'hc2f6b8cd;
    ram_cell[     187] = 32'h0;  // 32'h44873bc9;
    ram_cell[     188] = 32'h0;  // 32'h798458f7;
    ram_cell[     189] = 32'h0;  // 32'hb9a60f5c;
    ram_cell[     190] = 32'h0;  // 32'ha631ad8b;
    ram_cell[     191] = 32'h0;  // 32'h213d597a;
    ram_cell[     192] = 32'h0;  // 32'h75c5d6ea;
    ram_cell[     193] = 32'h0;  // 32'h2c308048;
    ram_cell[     194] = 32'h0;  // 32'h7265c120;
    ram_cell[     195] = 32'h0;  // 32'hd6fd4b51;
    ram_cell[     196] = 32'h0;  // 32'h60c12870;
    ram_cell[     197] = 32'h0;  // 32'h53663421;
    ram_cell[     198] = 32'h0;  // 32'h92cdab96;
    ram_cell[     199] = 32'h0;  // 32'h14bb647e;
    ram_cell[     200] = 32'h0;  // 32'hcadb8ff3;
    ram_cell[     201] = 32'h0;  // 32'hd7243f52;
    ram_cell[     202] = 32'h0;  // 32'ha9d3c39f;
    ram_cell[     203] = 32'h0;  // 32'h7398154c;
    ram_cell[     204] = 32'h0;  // 32'h0ee6982c;
    ram_cell[     205] = 32'h0;  // 32'h8fc2bf16;
    ram_cell[     206] = 32'h0;  // 32'hb4bd9fab;
    ram_cell[     207] = 32'h0;  // 32'h4887c468;
    ram_cell[     208] = 32'h0;  // 32'hd3e9a753;
    ram_cell[     209] = 32'h0;  // 32'hd68cee72;
    ram_cell[     210] = 32'h0;  // 32'h7f5470f4;
    ram_cell[     211] = 32'h0;  // 32'hb4bb8910;
    ram_cell[     212] = 32'h0;  // 32'h695eea78;
    ram_cell[     213] = 32'h0;  // 32'h815e3347;
    ram_cell[     214] = 32'h0;  // 32'h6f6a7e2a;
    ram_cell[     215] = 32'h0;  // 32'h9b9ea86a;
    ram_cell[     216] = 32'h0;  // 32'he2f3ad7b;
    ram_cell[     217] = 32'h0;  // 32'he66a5c22;
    ram_cell[     218] = 32'h0;  // 32'hd8a2b119;
    ram_cell[     219] = 32'h0;  // 32'ha3b4c918;
    ram_cell[     220] = 32'h0;  // 32'h83288610;
    ram_cell[     221] = 32'h0;  // 32'h755b1819;
    ram_cell[     222] = 32'h0;  // 32'h673c28aa;
    ram_cell[     223] = 32'h0;  // 32'he2451bc1;
    ram_cell[     224] = 32'h0;  // 32'h5d680c4e;
    ram_cell[     225] = 32'h0;  // 32'h8bbccc55;
    ram_cell[     226] = 32'h0;  // 32'h2efcd3be;
    ram_cell[     227] = 32'h0;  // 32'h902af0c9;
    ram_cell[     228] = 32'h0;  // 32'hfd6cf3b6;
    ram_cell[     229] = 32'h0;  // 32'h2f094ba2;
    ram_cell[     230] = 32'h0;  // 32'hab1eeea0;
    ram_cell[     231] = 32'h0;  // 32'h008286df;
    ram_cell[     232] = 32'h0;  // 32'hb687c82c;
    ram_cell[     233] = 32'h0;  // 32'h5ff5cc2c;
    ram_cell[     234] = 32'h0;  // 32'h7ebfe167;
    ram_cell[     235] = 32'h0;  // 32'h90f6a1e8;
    ram_cell[     236] = 32'h0;  // 32'h1ae82cb6;
    ram_cell[     237] = 32'h0;  // 32'h86896f87;
    ram_cell[     238] = 32'h0;  // 32'h583f29fc;
    ram_cell[     239] = 32'h0;  // 32'h69e3c0a5;
    ram_cell[     240] = 32'h0;  // 32'h907f325f;
    ram_cell[     241] = 32'h0;  // 32'hc1d68731;
    ram_cell[     242] = 32'h0;  // 32'hfb12e3c4;
    ram_cell[     243] = 32'h0;  // 32'ha3816dc3;
    ram_cell[     244] = 32'h0;  // 32'h7e70b1a2;
    ram_cell[     245] = 32'h0;  // 32'hc1272236;
    ram_cell[     246] = 32'h0;  // 32'h41326c25;
    ram_cell[     247] = 32'h0;  // 32'h88282a79;
    ram_cell[     248] = 32'h0;  // 32'ha588cf9d;
    ram_cell[     249] = 32'h0;  // 32'h9910abd5;
    ram_cell[     250] = 32'h0;  // 32'h274fc340;
    ram_cell[     251] = 32'h0;  // 32'h0020c559;
    ram_cell[     252] = 32'h0;  // 32'hd624b524;
    ram_cell[     253] = 32'h0;  // 32'h2a9ac5f6;
    ram_cell[     254] = 32'h0;  // 32'h9eb5dc1d;
    ram_cell[     255] = 32'h0;  // 32'h57ef58e8;
    // src matrix A
    ram_cell[     256] = 32'h3f2cb8c0;
    ram_cell[     257] = 32'h6972a8a4;
    ram_cell[     258] = 32'h15710b86;
    ram_cell[     259] = 32'h8085fdfc;
    ram_cell[     260] = 32'h25857d3d;
    ram_cell[     261] = 32'hd321337a;
    ram_cell[     262] = 32'he38e7d1b;
    ram_cell[     263] = 32'h56165f8c;
    ram_cell[     264] = 32'h8c7b6c9d;
    ram_cell[     265] = 32'hbfabe9b6;
    ram_cell[     266] = 32'h588aaa5b;
    ram_cell[     267] = 32'hb8b9e1d0;
    ram_cell[     268] = 32'hc96db5d6;
    ram_cell[     269] = 32'h7b136699;
    ram_cell[     270] = 32'h9c54edfa;
    ram_cell[     271] = 32'h15f256eb;
    ram_cell[     272] = 32'hfb3bb181;
    ram_cell[     273] = 32'h5bf80354;
    ram_cell[     274] = 32'he228386b;
    ram_cell[     275] = 32'hae882e9b;
    ram_cell[     276] = 32'h3c1fd1a0;
    ram_cell[     277] = 32'hb340dd6d;
    ram_cell[     278] = 32'hf310faeb;
    ram_cell[     279] = 32'h9556cf3d;
    ram_cell[     280] = 32'h6c16456b;
    ram_cell[     281] = 32'h50e3a0e5;
    ram_cell[     282] = 32'h14293cef;
    ram_cell[     283] = 32'he9ca4b00;
    ram_cell[     284] = 32'h04704a48;
    ram_cell[     285] = 32'h28611963;
    ram_cell[     286] = 32'h8c36d389;
    ram_cell[     287] = 32'h6ed56ca1;
    ram_cell[     288] = 32'h7a272a7b;
    ram_cell[     289] = 32'ha8a793e7;
    ram_cell[     290] = 32'hfb2ad2a5;
    ram_cell[     291] = 32'h5eec6efa;
    ram_cell[     292] = 32'h026b7c46;
    ram_cell[     293] = 32'h344c207f;
    ram_cell[     294] = 32'h3fb7ee57;
    ram_cell[     295] = 32'h0ab5ace0;
    ram_cell[     296] = 32'h7df22da1;
    ram_cell[     297] = 32'h7c31d5a0;
    ram_cell[     298] = 32'hbef9f622;
    ram_cell[     299] = 32'h6d1c587d;
    ram_cell[     300] = 32'h63290870;
    ram_cell[     301] = 32'h44469fa1;
    ram_cell[     302] = 32'hd15d9428;
    ram_cell[     303] = 32'h7ec787e3;
    ram_cell[     304] = 32'h9f48b3d8;
    ram_cell[     305] = 32'h40e3bdda;
    ram_cell[     306] = 32'h0f748ec6;
    ram_cell[     307] = 32'h47cbb2c9;
    ram_cell[     308] = 32'hf18b9d57;
    ram_cell[     309] = 32'h59eaecbe;
    ram_cell[     310] = 32'ha54cb7ef;
    ram_cell[     311] = 32'h0cc0a955;
    ram_cell[     312] = 32'he5fbd95f;
    ram_cell[     313] = 32'h9e64e100;
    ram_cell[     314] = 32'hd2c1b4eb;
    ram_cell[     315] = 32'hb43c3fdb;
    ram_cell[     316] = 32'hb95638e4;
    ram_cell[     317] = 32'ha10c8af4;
    ram_cell[     318] = 32'h103de0f5;
    ram_cell[     319] = 32'h7a3e9c20;
    ram_cell[     320] = 32'h302535a7;
    ram_cell[     321] = 32'h57c88423;
    ram_cell[     322] = 32'he6031ac1;
    ram_cell[     323] = 32'h7aaddd52;
    ram_cell[     324] = 32'h5538c7f5;
    ram_cell[     325] = 32'ha2968a7c;
    ram_cell[     326] = 32'hab132064;
    ram_cell[     327] = 32'h7d4436cb;
    ram_cell[     328] = 32'h975be63e;
    ram_cell[     329] = 32'ha2814e2b;
    ram_cell[     330] = 32'h90bb4b77;
    ram_cell[     331] = 32'he62eddac;
    ram_cell[     332] = 32'h41c81d5d;
    ram_cell[     333] = 32'hff8aa3c4;
    ram_cell[     334] = 32'h766e1d35;
    ram_cell[     335] = 32'h9f842d68;
    ram_cell[     336] = 32'h6dd35477;
    ram_cell[     337] = 32'h12a3633f;
    ram_cell[     338] = 32'hd3d2d2e3;
    ram_cell[     339] = 32'hdfa4364f;
    ram_cell[     340] = 32'he66fc760;
    ram_cell[     341] = 32'h12ed9f3d;
    ram_cell[     342] = 32'hdf20e523;
    ram_cell[     343] = 32'h55b16e73;
    ram_cell[     344] = 32'hdf202bc5;
    ram_cell[     345] = 32'h67e1e900;
    ram_cell[     346] = 32'hfb788639;
    ram_cell[     347] = 32'haeecd22d;
    ram_cell[     348] = 32'hec8bf7e3;
    ram_cell[     349] = 32'h58439efd;
    ram_cell[     350] = 32'h9d61b9c0;
    ram_cell[     351] = 32'hb12bac3f;
    ram_cell[     352] = 32'ha86b7e54;
    ram_cell[     353] = 32'h6e92b6c5;
    ram_cell[     354] = 32'h80481169;
    ram_cell[     355] = 32'h7e4ff882;
    ram_cell[     356] = 32'h3f2ecd03;
    ram_cell[     357] = 32'hf97041e8;
    ram_cell[     358] = 32'hdd96443b;
    ram_cell[     359] = 32'h2a93de77;
    ram_cell[     360] = 32'h1b11f11a;
    ram_cell[     361] = 32'h4786dede;
    ram_cell[     362] = 32'h11406db7;
    ram_cell[     363] = 32'ha7a5347c;
    ram_cell[     364] = 32'hb60e2348;
    ram_cell[     365] = 32'h3d252029;
    ram_cell[     366] = 32'h1c19db1c;
    ram_cell[     367] = 32'hbfc88283;
    ram_cell[     368] = 32'h997287cb;
    ram_cell[     369] = 32'h91d95014;
    ram_cell[     370] = 32'hc3f31997;
    ram_cell[     371] = 32'hddc072dc;
    ram_cell[     372] = 32'h6a579270;
    ram_cell[     373] = 32'h1a53e246;
    ram_cell[     374] = 32'hd33fc155;
    ram_cell[     375] = 32'h8e329396;
    ram_cell[     376] = 32'h0c16531d;
    ram_cell[     377] = 32'hf7a8282d;
    ram_cell[     378] = 32'h3eef2777;
    ram_cell[     379] = 32'h4e42647a;
    ram_cell[     380] = 32'habe39d50;
    ram_cell[     381] = 32'h1d7cf35d;
    ram_cell[     382] = 32'hdbb8821b;
    ram_cell[     383] = 32'hd46cd5a8;
    ram_cell[     384] = 32'h5aefac2d;
    ram_cell[     385] = 32'hbb28b1a3;
    ram_cell[     386] = 32'h2c378567;
    ram_cell[     387] = 32'he3a910bb;
    ram_cell[     388] = 32'hea25a5a6;
    ram_cell[     389] = 32'hcff56036;
    ram_cell[     390] = 32'h1d6b82c9;
    ram_cell[     391] = 32'h90c24c54;
    ram_cell[     392] = 32'h45999cfa;
    ram_cell[     393] = 32'heca77f33;
    ram_cell[     394] = 32'hbfe97bfd;
    ram_cell[     395] = 32'hbbcdb65e;
    ram_cell[     396] = 32'hbc26b8a2;
    ram_cell[     397] = 32'h8291e062;
    ram_cell[     398] = 32'hc4302de0;
    ram_cell[     399] = 32'hd8ac84f3;
    ram_cell[     400] = 32'hc9bb0b35;
    ram_cell[     401] = 32'h861e2183;
    ram_cell[     402] = 32'h6747f283;
    ram_cell[     403] = 32'h1bdbe5ae;
    ram_cell[     404] = 32'hf5000aa2;
    ram_cell[     405] = 32'h6bd2a446;
    ram_cell[     406] = 32'hecb06d06;
    ram_cell[     407] = 32'hd9e3d899;
    ram_cell[     408] = 32'h70818d20;
    ram_cell[     409] = 32'h0c8a8c69;
    ram_cell[     410] = 32'hceff3ac6;
    ram_cell[     411] = 32'h1b4bc289;
    ram_cell[     412] = 32'hc515e723;
    ram_cell[     413] = 32'h5ac9487a;
    ram_cell[     414] = 32'h12717968;
    ram_cell[     415] = 32'had39ee31;
    ram_cell[     416] = 32'h6e6bcc18;
    ram_cell[     417] = 32'h8104868f;
    ram_cell[     418] = 32'hb3d74510;
    ram_cell[     419] = 32'h2bb8fd9f;
    ram_cell[     420] = 32'hc2108ff6;
    ram_cell[     421] = 32'h4fa2ec3a;
    ram_cell[     422] = 32'h29d2aa55;
    ram_cell[     423] = 32'hf6f1eaaf;
    ram_cell[     424] = 32'h0a3d085d;
    ram_cell[     425] = 32'h1b85ebf6;
    ram_cell[     426] = 32'h8dad2587;
    ram_cell[     427] = 32'hcfdf14e3;
    ram_cell[     428] = 32'h4e1eae2b;
    ram_cell[     429] = 32'hfb6cda7e;
    ram_cell[     430] = 32'h804fb6b7;
    ram_cell[     431] = 32'h2b824a6a;
    ram_cell[     432] = 32'h69341508;
    ram_cell[     433] = 32'h554396e4;
    ram_cell[     434] = 32'h35ea48f8;
    ram_cell[     435] = 32'h5518ed2a;
    ram_cell[     436] = 32'hd30f5963;
    ram_cell[     437] = 32'h8db7873e;
    ram_cell[     438] = 32'h6417b5e7;
    ram_cell[     439] = 32'h0da8df0f;
    ram_cell[     440] = 32'hae75c7e0;
    ram_cell[     441] = 32'hbdfef117;
    ram_cell[     442] = 32'h19b0d979;
    ram_cell[     443] = 32'hc9bbde9a;
    ram_cell[     444] = 32'h409cdf17;
    ram_cell[     445] = 32'h2f78001c;
    ram_cell[     446] = 32'h9349c465;
    ram_cell[     447] = 32'hbf6222ec;
    ram_cell[     448] = 32'h2b866566;
    ram_cell[     449] = 32'h08623f90;
    ram_cell[     450] = 32'h1bbe17cc;
    ram_cell[     451] = 32'h43bb267b;
    ram_cell[     452] = 32'h973e22cb;
    ram_cell[     453] = 32'hebc1eae3;
    ram_cell[     454] = 32'h3fc62778;
    ram_cell[     455] = 32'h58a5b72f;
    ram_cell[     456] = 32'h30958149;
    ram_cell[     457] = 32'ha9023c2e;
    ram_cell[     458] = 32'h593df3a7;
    ram_cell[     459] = 32'ha4330014;
    ram_cell[     460] = 32'h5dd2e055;
    ram_cell[     461] = 32'h8a18381c;
    ram_cell[     462] = 32'h5cae2f31;
    ram_cell[     463] = 32'h22954203;
    ram_cell[     464] = 32'hd2aa7f71;
    ram_cell[     465] = 32'h17e10e78;
    ram_cell[     466] = 32'hd6c1e834;
    ram_cell[     467] = 32'hb8306d35;
    ram_cell[     468] = 32'h5e5be526;
    ram_cell[     469] = 32'hc2e62b4b;
    ram_cell[     470] = 32'h37a0ad1c;
    ram_cell[     471] = 32'hc56c3cf3;
    ram_cell[     472] = 32'h98003c0e;
    ram_cell[     473] = 32'h3a968066;
    ram_cell[     474] = 32'h2aabc7f6;
    ram_cell[     475] = 32'hcd0bdb5d;
    ram_cell[     476] = 32'h56d9dc29;
    ram_cell[     477] = 32'h179f8089;
    ram_cell[     478] = 32'hca711582;
    ram_cell[     479] = 32'h535eb60c;
    ram_cell[     480] = 32'h2b373548;
    ram_cell[     481] = 32'h088c73ac;
    ram_cell[     482] = 32'h328a8d4d;
    ram_cell[     483] = 32'h2e4597c9;
    ram_cell[     484] = 32'h032419df;
    ram_cell[     485] = 32'h45267d05;
    ram_cell[     486] = 32'hdcbb6716;
    ram_cell[     487] = 32'h01430326;
    ram_cell[     488] = 32'h3d64120b;
    ram_cell[     489] = 32'h08fecd45;
    ram_cell[     490] = 32'h4e66a82b;
    ram_cell[     491] = 32'h66eaa136;
    ram_cell[     492] = 32'h8dcb879d;
    ram_cell[     493] = 32'h7b5a4cdc;
    ram_cell[     494] = 32'hacfb41b6;
    ram_cell[     495] = 32'hdb2587a4;
    ram_cell[     496] = 32'hf1e0b233;
    ram_cell[     497] = 32'hfebd46b0;
    ram_cell[     498] = 32'hd11f7f81;
    ram_cell[     499] = 32'h135f45e2;
    ram_cell[     500] = 32'h92b5fac5;
    ram_cell[     501] = 32'h4f97b6f3;
    ram_cell[     502] = 32'h578d569e;
    ram_cell[     503] = 32'hfdd6b4d3;
    ram_cell[     504] = 32'h0584be9d;
    ram_cell[     505] = 32'hf8150fc1;
    ram_cell[     506] = 32'hae1a9abc;
    ram_cell[     507] = 32'h2bf17378;
    ram_cell[     508] = 32'h3d6ceba9;
    ram_cell[     509] = 32'h2d83abb4;
    ram_cell[     510] = 32'h71fca7e1;
    ram_cell[     511] = 32'h614cc785;
    // src matrix B
    ram_cell[     512] = 32'hb3a89d70;
    ram_cell[     513] = 32'h8e56ceaf;
    ram_cell[     514] = 32'h4546779c;
    ram_cell[     515] = 32'h8f4db8d5;
    ram_cell[     516] = 32'h43b455af;
    ram_cell[     517] = 32'h628daa0d;
    ram_cell[     518] = 32'hb6460e93;
    ram_cell[     519] = 32'he13b5c41;
    ram_cell[     520] = 32'hfd6f4089;
    ram_cell[     521] = 32'hba78ef35;
    ram_cell[     522] = 32'h397fb892;
    ram_cell[     523] = 32'hd2379e54;
    ram_cell[     524] = 32'h377d25ec;
    ram_cell[     525] = 32'hcd3d5713;
    ram_cell[     526] = 32'hd1b7c2e3;
    ram_cell[     527] = 32'hed247415;
    ram_cell[     528] = 32'h4baca4c8;
    ram_cell[     529] = 32'h094a536b;
    ram_cell[     530] = 32'h2406f195;
    ram_cell[     531] = 32'h815f1ed4;
    ram_cell[     532] = 32'he0ae6b90;
    ram_cell[     533] = 32'hfed0e35d;
    ram_cell[     534] = 32'he89635bb;
    ram_cell[     535] = 32'h9b083ab1;
    ram_cell[     536] = 32'h6280d820;
    ram_cell[     537] = 32'h837e273c;
    ram_cell[     538] = 32'h1f13cf88;
    ram_cell[     539] = 32'h9725a779;
    ram_cell[     540] = 32'h5a0134c6;
    ram_cell[     541] = 32'hef512f36;
    ram_cell[     542] = 32'h1ee037d9;
    ram_cell[     543] = 32'hf7771207;
    ram_cell[     544] = 32'h8a7cce54;
    ram_cell[     545] = 32'h3813978a;
    ram_cell[     546] = 32'h0821b402;
    ram_cell[     547] = 32'h4be372d4;
    ram_cell[     548] = 32'h6ef94311;
    ram_cell[     549] = 32'h3e88e382;
    ram_cell[     550] = 32'h1fb05acc;
    ram_cell[     551] = 32'h47dfe0bd;
    ram_cell[     552] = 32'heeae33ef;
    ram_cell[     553] = 32'h298ae1b3;
    ram_cell[     554] = 32'h726606e2;
    ram_cell[     555] = 32'hd3da65c9;
    ram_cell[     556] = 32'h3de5f282;
    ram_cell[     557] = 32'hdb044b0e;
    ram_cell[     558] = 32'h7794a544;
    ram_cell[     559] = 32'hc2738860;
    ram_cell[     560] = 32'h9c06561a;
    ram_cell[     561] = 32'h14cbb19d;
    ram_cell[     562] = 32'h41803573;
    ram_cell[     563] = 32'h12e7ff2c;
    ram_cell[     564] = 32'he7ce60be;
    ram_cell[     565] = 32'h44928e37;
    ram_cell[     566] = 32'h3452929c;
    ram_cell[     567] = 32'h067f4d42;
    ram_cell[     568] = 32'h8968d7d2;
    ram_cell[     569] = 32'h50ca1cd4;
    ram_cell[     570] = 32'h0bb94116;
    ram_cell[     571] = 32'hd2eaa10a;
    ram_cell[     572] = 32'h1d1a54fe;
    ram_cell[     573] = 32'hfc30e6eb;
    ram_cell[     574] = 32'he64be081;
    ram_cell[     575] = 32'h9db1c34c;
    ram_cell[     576] = 32'h1d9ec83e;
    ram_cell[     577] = 32'h8f1e3bba;
    ram_cell[     578] = 32'hb085a092;
    ram_cell[     579] = 32'hdfcab2f3;
    ram_cell[     580] = 32'hb338429e;
    ram_cell[     581] = 32'hf230a562;
    ram_cell[     582] = 32'h1e3ebeff;
    ram_cell[     583] = 32'h87f6af10;
    ram_cell[     584] = 32'hf429b7da;
    ram_cell[     585] = 32'hea9000b9;
    ram_cell[     586] = 32'h48614cc1;
    ram_cell[     587] = 32'h8d5b9fa2;
    ram_cell[     588] = 32'hf360b66a;
    ram_cell[     589] = 32'h3a3f4f2d;
    ram_cell[     590] = 32'h574c065b;
    ram_cell[     591] = 32'heae5a7d7;
    ram_cell[     592] = 32'hd6211952;
    ram_cell[     593] = 32'h8465a522;
    ram_cell[     594] = 32'h983a0483;
    ram_cell[     595] = 32'h3c659b91;
    ram_cell[     596] = 32'hc66f2c2f;
    ram_cell[     597] = 32'h80c89f1a;
    ram_cell[     598] = 32'hc2966329;
    ram_cell[     599] = 32'h34bfbc67;
    ram_cell[     600] = 32'h0879cede;
    ram_cell[     601] = 32'hab92f7aa;
    ram_cell[     602] = 32'h15e6fd1f;
    ram_cell[     603] = 32'h67e71025;
    ram_cell[     604] = 32'hc53c14ff;
    ram_cell[     605] = 32'hb451c284;
    ram_cell[     606] = 32'h883cae12;
    ram_cell[     607] = 32'hf5a42cba;
    ram_cell[     608] = 32'hf6aede28;
    ram_cell[     609] = 32'hcc48f8f0;
    ram_cell[     610] = 32'h380d08ea;
    ram_cell[     611] = 32'hb1b90b7d;
    ram_cell[     612] = 32'ha8288b85;
    ram_cell[     613] = 32'h67656a85;
    ram_cell[     614] = 32'h084bb548;
    ram_cell[     615] = 32'h29e571b1;
    ram_cell[     616] = 32'hd8665d85;
    ram_cell[     617] = 32'h0ae60935;
    ram_cell[     618] = 32'h33ed0a9a;
    ram_cell[     619] = 32'hf2a0356b;
    ram_cell[     620] = 32'h57735c0b;
    ram_cell[     621] = 32'h1f5e6a4c;
    ram_cell[     622] = 32'h33d5f2d5;
    ram_cell[     623] = 32'hed7badde;
    ram_cell[     624] = 32'ha810195f;
    ram_cell[     625] = 32'hf9068715;
    ram_cell[     626] = 32'h8c101ea2;
    ram_cell[     627] = 32'h40cc7b5b;
    ram_cell[     628] = 32'h808e624e;
    ram_cell[     629] = 32'hb4e2ae39;
    ram_cell[     630] = 32'hf3f587bf;
    ram_cell[     631] = 32'h1069632d;
    ram_cell[     632] = 32'h7679eb75;
    ram_cell[     633] = 32'h936a845e;
    ram_cell[     634] = 32'hfbd1e711;
    ram_cell[     635] = 32'h27159f71;
    ram_cell[     636] = 32'hcc45be75;
    ram_cell[     637] = 32'ha54e4e80;
    ram_cell[     638] = 32'hccfb1713;
    ram_cell[     639] = 32'ha77dd3b1;
    ram_cell[     640] = 32'h153996fe;
    ram_cell[     641] = 32'hae3e83c1;
    ram_cell[     642] = 32'hfcadcbd5;
    ram_cell[     643] = 32'h6c58c502;
    ram_cell[     644] = 32'hf45b9c23;
    ram_cell[     645] = 32'h9f285fdb;
    ram_cell[     646] = 32'h853a2ea6;
    ram_cell[     647] = 32'hec59287b;
    ram_cell[     648] = 32'h8430acfb;
    ram_cell[     649] = 32'hf54d6f2f;
    ram_cell[     650] = 32'h26570f64;
    ram_cell[     651] = 32'h276b1ff2;
    ram_cell[     652] = 32'ha25eea37;
    ram_cell[     653] = 32'hca6d7873;
    ram_cell[     654] = 32'hcc254e3c;
    ram_cell[     655] = 32'h2459af48;
    ram_cell[     656] = 32'he84d42e5;
    ram_cell[     657] = 32'h40254f29;
    ram_cell[     658] = 32'hae30dc28;
    ram_cell[     659] = 32'hcd60ce1b;
    ram_cell[     660] = 32'h391569d6;
    ram_cell[     661] = 32'hd20241af;
    ram_cell[     662] = 32'h366618cf;
    ram_cell[     663] = 32'h856ba197;
    ram_cell[     664] = 32'h9f66fed0;
    ram_cell[     665] = 32'h576280bf;
    ram_cell[     666] = 32'ha947878d;
    ram_cell[     667] = 32'heb4aa8e0;
    ram_cell[     668] = 32'h32457035;
    ram_cell[     669] = 32'hf0ced407;
    ram_cell[     670] = 32'h7cd354d6;
    ram_cell[     671] = 32'h55a84370;
    ram_cell[     672] = 32'h5a52b5d8;
    ram_cell[     673] = 32'had1e21b6;
    ram_cell[     674] = 32'h2a3dd8d5;
    ram_cell[     675] = 32'hc6e9bb32;
    ram_cell[     676] = 32'h7a55c7bc;
    ram_cell[     677] = 32'hd7912870;
    ram_cell[     678] = 32'h3c22bd83;
    ram_cell[     679] = 32'hacaa55ae;
    ram_cell[     680] = 32'h7d65b586;
    ram_cell[     681] = 32'h383258dc;
    ram_cell[     682] = 32'hf6210340;
    ram_cell[     683] = 32'h5210483e;
    ram_cell[     684] = 32'h6cf60eb9;
    ram_cell[     685] = 32'h003b1237;
    ram_cell[     686] = 32'h5ba9cca8;
    ram_cell[     687] = 32'ha1ced56b;
    ram_cell[     688] = 32'h1960c973;
    ram_cell[     689] = 32'h572916be;
    ram_cell[     690] = 32'hcda4fcdc;
    ram_cell[     691] = 32'hfea2ae50;
    ram_cell[     692] = 32'h973ee09f;
    ram_cell[     693] = 32'h0e5bc435;
    ram_cell[     694] = 32'ha015d2fd;
    ram_cell[     695] = 32'h7f85042b;
    ram_cell[     696] = 32'ha9f79508;
    ram_cell[     697] = 32'ha8bd3d6c;
    ram_cell[     698] = 32'h3bdb5feb;
    ram_cell[     699] = 32'hcf36b41a;
    ram_cell[     700] = 32'h730fc34b;
    ram_cell[     701] = 32'hfca9389f;
    ram_cell[     702] = 32'ha0fb8a49;
    ram_cell[     703] = 32'he19fced8;
    ram_cell[     704] = 32'hdcc22ea7;
    ram_cell[     705] = 32'h1a65428c;
    ram_cell[     706] = 32'h7d9e1ae6;
    ram_cell[     707] = 32'h1e2d7e58;
    ram_cell[     708] = 32'h036c970f;
    ram_cell[     709] = 32'h86e50a31;
    ram_cell[     710] = 32'h67392ab0;
    ram_cell[     711] = 32'h667f2683;
    ram_cell[     712] = 32'h8016f6de;
    ram_cell[     713] = 32'ha618b30c;
    ram_cell[     714] = 32'h156e8392;
    ram_cell[     715] = 32'hef5e6bc2;
    ram_cell[     716] = 32'h74419328;
    ram_cell[     717] = 32'hf6a9b1a2;
    ram_cell[     718] = 32'hcc4bf904;
    ram_cell[     719] = 32'h6f7e7fc5;
    ram_cell[     720] = 32'hb2e8a9f6;
    ram_cell[     721] = 32'h5b45b7d9;
    ram_cell[     722] = 32'h10ae6df0;
    ram_cell[     723] = 32'h969b075d;
    ram_cell[     724] = 32'h463fd7c2;
    ram_cell[     725] = 32'hd99913a0;
    ram_cell[     726] = 32'h9bc74108;
    ram_cell[     727] = 32'hd04f454b;
    ram_cell[     728] = 32'h403e7121;
    ram_cell[     729] = 32'h7b2a5513;
    ram_cell[     730] = 32'h7e54af80;
    ram_cell[     731] = 32'h6da4f4f0;
    ram_cell[     732] = 32'h495bd75f;
    ram_cell[     733] = 32'hf8834028;
    ram_cell[     734] = 32'hde711b42;
    ram_cell[     735] = 32'h6a08e86c;
    ram_cell[     736] = 32'h9ba3d5d5;
    ram_cell[     737] = 32'hc614762d;
    ram_cell[     738] = 32'h8df7e279;
    ram_cell[     739] = 32'he2684d2a;
    ram_cell[     740] = 32'h5a299946;
    ram_cell[     741] = 32'h9235437a;
    ram_cell[     742] = 32'h74481084;
    ram_cell[     743] = 32'hd26d50a5;
    ram_cell[     744] = 32'h8e820ac5;
    ram_cell[     745] = 32'ha260119c;
    ram_cell[     746] = 32'h5f25cbd0;
    ram_cell[     747] = 32'haef519d5;
    ram_cell[     748] = 32'hb2c5575f;
    ram_cell[     749] = 32'h314efeb1;
    ram_cell[     750] = 32'he20f9ea2;
    ram_cell[     751] = 32'hf1e33d9c;
    ram_cell[     752] = 32'h7eb40fb3;
    ram_cell[     753] = 32'h0f78661c;
    ram_cell[     754] = 32'hd8fb37f3;
    ram_cell[     755] = 32'h68c5d70e;
    ram_cell[     756] = 32'h092959e9;
    ram_cell[     757] = 32'hc09a7011;
    ram_cell[     758] = 32'ha86956dc;
    ram_cell[     759] = 32'h6e8a44a9;
    ram_cell[     760] = 32'hc35d8494;
    ram_cell[     761] = 32'h2ab76bfa;
    ram_cell[     762] = 32'hf96ee40a;
    ram_cell[     763] = 32'h09f91677;
    ram_cell[     764] = 32'h5db43401;
    ram_cell[     765] = 32'ha9925441;
    ram_cell[     766] = 32'hdb61fee6;
    ram_cell[     767] = 32'ha406ec76;
end

endmodule

